/********************************************************
# Description: definition of the hard adder black-box	#
#														#
# Author: Seyed Alireza Damghani (sdamghann@gmail.com)  #
********************************************************/

(* blackbox *)
module adder(a, b, cin, cout, sumout);
	input a, b, cin;
	output cout, sumout;
	
	//assign {cout,sumout} = a + b + cin;
endmodule
